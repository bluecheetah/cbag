*.BIPOLAR
*.RESI = 2000
*.SCALE METER
*.MEGA
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
.PARAM


.SUBCKT TEST B D G S
*.PININFO B:B D:B G:B S:B
.ENDS
