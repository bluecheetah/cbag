*.BIPOLAR
*.RESI = 2000
*.SCALE METER
*.MEGA
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
.PARAM


.SUBCKT pmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
.ENDS


.SUBCKT TEST VDD VSS in out
*.PININFO VDD:I VSS:I in:I out:O
XP VDD out in VSS / pmos4_standard l=90n nf=2 w=400n
.ENDS
