*.BIPOLAR
*.RESI = 2000
*.SCALE METER
*.MEGA
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
.PARAM


.SUBCKT pmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
.ENDS


.SUBCKT cv_bus_term VDD VSS in<1> in<0> out
*.PININFO VDD:I VSS:I in<1>:I in<0>:I out:O
X4 VDD out in<1> VSS / pmos4_standard l=90n nf=2 w=400n
XP VDD out in<0> VSS / pmos4_standard l=90n nf=2 w=400n
.ENDS


.SUBCKT TEST VDD VSS in<1> in<0> out
*.PININFO VDD:I VSS:I in<1>:I in<0>:I out:O
XINST VDD VSS in<1> in<0> out / cv_bus_term
.ENDS
