*.BIPOLAR
*.RESI = 2000
*.SCALE METER
*.MEGA
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
.PARAM


.SUBCKT nmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
.ENDS


.SUBCKT pmos4_standard B D G S
*.PININFO B:B D:B G:B S:B
.ENDS


.SUBCKT TEST VDD VSS in out
*.PININFO VDD:I VSS:I in:I out:O
XN VSS out in VSS / nmos4_standard
XP VDD out in VDD / pmos4_standard l=90n nf=2 w=400n
.ENDS
