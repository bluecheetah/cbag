

module TEST(
    input  wire VDD,
    input  wire VSS,
    input  wire [1:0] in0,
    input  wire [1:0] in1,
    output wire [1:0] out
);

endmodule
